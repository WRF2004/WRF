module comparator (
	input[3:0] A,    
	input[3:0] B, 
	output Out
);
wire[3:0] a;
wire[3:0] b;
assign a = ~A + 1;
assign b = ~B + 1;
assign Out = (A[3] == 1 && B[3] == 0) ? 1 : (A[3] == 0 && B[3] == 1) ? 0 :
			 ((A[3] == 0 && B[3] == 0) && (A[2] == 0 && B[2] == 1)) ? 1 :
			 ((A[3] == 0 && B[3] == 0) && (A[2] == 1 && B[2] == 0)) ? 0 :
			 ((A[3] == 0 && B[3] == 0) && (A[1] == 0 && B[1] == 1)) ? 1 :
			 ((A[3] == 0 && B[3] == 0) && (A[1] == 1 && B[1] == 0)) ? 0 :
			 ((A[3] == 0 && B[3] == 0) && (A[0] == 0 && B[0] == 1)) ? 1 :
			 ((A[3] == 0 && B[3] == 0) && (A[0] == 1 && B[0] == 0)) ? 0 :
			 ((a[3] == 0 && b[3] == 0) && (a[2] == 1 && b[2] == 0)) ? 1 :
			 ((a[3] == 0 && b[3] == 0) && (a[2] == 0 && b[2] == 1)) ? 0 :
			 ((a[3] == 0 && b[3] == 0) && (a[1] == 1 && b[1] == 0)) ? 1 :
			 ((a[3] == 0 && b[3] == 0) && (a[1] == 0 && b[1] == 1)) ? 0 :
			 ((a[3] == 0 && b[3] == 0) && (a[0] == 1 && b[0] == 0)) ? 1 :
			 ((a[3] == 0 && b[3] == 0) && (a[0] == 0 && b[0] == 1)) ? 0 :
			 							(a[3] == 1 && b[3] == 0) ? 1 : 0; 

endmodule